module TriangularWave(input clk,output reg [15:0]Triangularout,input reset,input[6:0]phase);
endmodule
