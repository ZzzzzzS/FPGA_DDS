module ClockGenerator(input clk,input [1:0]Switch,input [1:0]SwitchMicro,input [1:0]SwitchNano,output reg clk_N,input reset);

endmodule
