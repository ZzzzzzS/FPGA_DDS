module phase (input add,input sub,output [6:0]phase,input reset);
endmodule
