module SinWave(input clk,output reg [15:0]Sinout,input reset,input[7:0]phase);
endmodule
