module PWMWave(input clk,input [7:0]PWMDuty,output reg [15:0]PWMout,input reset,input[6:0]phase);
endmodule
