module TriangularWave(input clk,output [15:0]Triangularout,input reset,input[31:0]phase,input[31:0]Step);
reg [31:0]address;
reg [31:0]SynthesisedPhase;
initial
    begin
        address=32'd0;
    end

TriangularROM ROM1(.address(SynthesisedPhase),
             .clock(clk),
             .q(Triangularout));

always@(negedge clk)
    begin
        address<=address+Step;
        SynthesisedPhase<=address+phase;
    end
endmodule
