module phase (input add,input sub,output [7:0]phase,input reset);
endmodule
